---Half Adder wrap---------
---library description-----
Library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--port description-----
entity half_adder is 
port (
    a,b  : in  std_logic;
	  sum  : out std_logic;
	  carry: out std_logic
	  );
end half_adder;

--architecture description-----
architecture behavioural of half_adder is 
begin

sum   <= a xor b;  --xor gate 
carry <= a and b;  --and gate

end behavioural;

---Full adder wrap using two-half adder------
---Library description------
Library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

---port description------
entity full_adder is
port(
   a,b,ci  : in  std_logic;
	 s       : out std_logic;
	 cout    : out std_logic
	 );
end full_adder;

---architecture description------
architecture behavioral of full_adder is
---signal,constants,component instant etc... description------
signal s_sig        : std_logic;
signal c_sig,c_sig1 : std_logic;
--------------------------------------------------------------
begin

---Instantiation------
HA1: entity work.half_adder
port map(
    a     => a,
    b     => b,
	  sum   => s_sig, 
	  carry => c_sig
	  );
   
HA2: entity work.half_adder
port map(
    a     => s_sig,
    b     => ci,
	  sum   => s ,
	  carry => c_sig1
	  );

cout <= c_sig or c_sig1;   
end behavioral; 